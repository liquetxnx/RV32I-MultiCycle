

`include "defines.v"
module stage_ID(
    input clk,
    input rst,

    input wire [31:0] if_instr,

    input wire [4:0] wb_rd,
    input wire [31:0] wb_wd,
    input wire wb_regwrite,

    output wire id_a_sel,
    output wire id_b_sel,
    output wire [1:0] id_alu_op,
    output wire [1:0] id_pc_op,
    output wire id_regwrite,
    output wire id_memwrite,
    output wire [1:0] id_memtoreg,

    output wire [31:0] id_imm,
    output wire [3:0] id_funct3,
    output wire [4:0] id_rd,

    output wire [31:0] id_rdata1,
    output wire [31:0] id_rdata2
);

wire [2:0] immsrc;

Control_Unit ctrl_inst(

    .opcode(if_instr[6:0]),

    .a_sel(id_a_sel),
    .b_sel(id_b_sel),
    .alu_op(id_alu_op),
    .pc_op(id_pc_op),
    .regwrite(id_regwrite),
    .memwrite(id_memwrite),
    .memtoreg(id_memtoreg),
    .immsrc(immsrc)
);

ImmGen immgen_inst(
    .instr(if_instr[31:7]),
    .immsrc(immsrc),
    .imm(id_imm)

);


Reg_File reg_inst(
    .clk(clk),
    .rst(rst),
    .regwrite(wb_regwrite),
    .rs1(if_instr[19:15]),
    .rs2(if_instr[24:20]),
    .rd(wb_rd),
    .wd(wb_wd),
    .rdata1(id_rdata1),
    .rdata2(id_rdata2)
);
assign id_funct3 = if_instr[14:12];
assign id_rd = if_instr[11:7];

endmodule
